
library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity InstMem is
  generic (BitWidth: integer;
           InstructionWidth: integer);
  port ( address : in std_logic_vector(BitWidth-1 downto 0);
         data : out std_logic_vector(InstructionWidth-1 downto 0) );
end entity InstMem;

architecture behavioral of InstMem is
  
  type mem is array ( 0 to (2**BitWidth)-1) of std_logic_vector(InstructionWidth-1 downto 0);
  
  constant my_InstMem : mem := (
	 0 =>   "01111100000011",
	 1 =>   "01010000000000",
	 2 =>   "01111100000011",
	 3 =>   "01010000000101",
	 4 =>   "01001100000010",
	 5 =>   "01111100000001",
	 6 =>   "00010100001000",
	 7 =>   "01010000010100",
	 8 =>   "01111100000001",
	 9 =>   "00010100000100",
	 10 =>   "01010000011000",
	 11 =>   "01111100000001",
	 12 =>   "00010100000010",
	 13 =>   "01010000011100",
	 14 =>   "01111100000001",
	 15 =>   "00010100000001",
	 16 =>   "01010000100010",
	 17 =>   "01111100000001",
	 18 =>   "00010100000001",
	 19 =>   "01001100000000",
	 20 =>   "01111100000100",
	 21 =>   "00000100000010",
	 22 =>   "10000000000100",
	 23 =>   "01001100000000",
	 24 =>   "01111100000100",
	 25 =>   "00010000000010",
	 26 =>   "10000000000100",
	 27 =>   "01001100000000",
	 28 =>   "01111100000100",
	 29 =>   "10010000000001",
	 30 =>   "01111100000010",
	 31 =>   "00111000000000",
	 32 =>   "10000000000100",
	 33 =>   "01001100000000",
	 34 =>   "01111100000100",
	 35 =>   "10010000000001",
	 36 =>   "01111100000010",
	 37 =>   "00111100000000",
	 38 =>   "10000000000100",
	 39 =>   "01001100000000",
others => "00000000000000"
    );
    

begin
  
  data <= my_InstMem(to_integer(unsigned(address)));

  
end architecture behavioral;